module hexdriver (input [3:0] val, output logic [6:0] HEX);

	/* your code here */
	// 0 ---> 0000
	// 1 ---> 0001
	// 2 ---> 0010
	// 3 ---> 0011
	// 4 ---> 0100
	// 5 ---> 0101
	// 6 ---> 0110
	// 7 ---> 0111
	// 8 ---> 1000
	// 9 ---> 1001
	// 10 --> 1010 (A)
	// 11 --> 1011 (B)
	// 12 --> 1100 (C)
	// 13 --> 1101 (D)
	// 14 --> 1110 (E)
	// 15 --> 1111 (F)
	
	always_comb begin
		case (val)
			4'd0: HEX = 7'b100_0000;  // 0
			4'd1: HEX = 7'b111_1001;  // 1
			4'd2: HEX = 7'b010_0100;  // 2
			4'd3: HEX = 7'b011_0000;  // 3
			4'd4: HEX = 7'b001_1001;  // 4
			4'd5: HEX = 7'b001_0010;  // 5
			4'd6: HEX = 7'b000_0010;  // 6
			4'd7: HEX = 7'b111_1000;  // 7
			4'd8: HEX = 7'b000_0000;  // 8
			4'd9: HEX = 7'b001_1000;  // 9
			4'd10: HEX = 7'b000_1000;  // A
			4'd11: HEX = 7'b000_0011;  // b
			4'd12: HEX = 7'b100_0110;  // C
			4'd13: HEX = 7'b010_0001;  // d
			4'd14: HEX = 7'b000_0110;  // E
			4'd15: HEX = 7'b000_1110;  // F
			default: HEX = 7'b000_0000;  // off
		endcase
	end
endmodule
