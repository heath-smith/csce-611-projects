module hexdriver (input [3:0] val, output logic [6:0] HEX);

	/* your code here */
	// 0 ---> 0000
	// 1 ---> 0001
	// 2 ---> 0010
	// 3 ---> 0011
	// 4 ---> 0100
	// 5 ---> 0101
	// 6 ---> 0110
	// 7 ---> 0111
	// 8 ---> 1000
	// 9 ---> 1001
	// 10 --> 1010 (A)
	// 11 --> 1011 (B)
	// 12 --> 1100 (C)
	// 13 --> 1101 (D)
	// 14 --> 1110 (E)
	// 15 --> 1111 (F)
	
	always_comb
		case (val)
			4'd0: HEX = 7'b011_1111;  // 0
			4'd1: HEX = 7'b000_0110;  // 1
			4'd2: HEX = 7'b101_1011;  // 2
			4'd3: HEX = 7'b100_1111;  // 3
			4'd4: HEX = 7'b110_0110;  // 4
			4'd5: HEX = 7'b110_1101;  // 5
			4'd6: HEX = 7'b111_1101;  // 6
			4'd7: HEX = 7'b000_0111;  // 7
			4'd8: HEX = 7'b111_1111;  // 8
			4'd9: HEX = 7'b110_0111;  // 9
			4'd10: HEX = 7'b111_0111;  // A
			4'd11: HEX = 7'b111_1100;  // b
			4'd12: HEX = 7'b011_1001;  // C
			4'd13: HEX = 7'b101_1110;  // d
			4'd14: HEX = 7'b111_1001;  // E
			4'd15: HEX = 7'b111_0001;  // F
			default: HEX = 7'b000_0000;  // off
	end

endmodule
