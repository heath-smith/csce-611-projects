// controller unit
module controller(

);

    always_comb begin
        // set defaults here
        if () begin
            //
        end else begin
            //
        end
    end

endmodule